module top( input logic MAX10_CLK1_50, 
           input logic [9:0] SW,
           input logic [1:0] KEY,
    		output logic [31:0] WriteData, DataAdr,
    		output logic MemWrite,
           output logic [9:0] LEDR,
			  output logic [7:0] HEX0,
			  output logic [7:0] HEX1,
			  output logic [7:0] HEX2,
			  output logic [7:0] HEX3,
			  output logic [7:0] HEX4,
			  output logic [7:0] HEX5);

			logic clk;
			assign clk = MAX10_CLK1_50;
			
			logic [15:0] HEX5HEX4;
			logic [31:0] HEX3HEX0;
			
			assign {HEX3,HEX2,HEX1,HEX0} = ~HEX3HEX0;
			assign {HEX5,HEX4} = ~HEX5HEX4;
			
  logic [31:0] PC, Instr, ReadData, MemReadData;
  
  logic reset;
  assign reset = ~KEY[1];
  
    // instantiate processor and memories
  riscvsingle rvsingle(clk, reset, PC, Instr, MemWrite, DataAdr,	  WriteData, ReadData);
  imem imem(PC, Instr);
  dmem dmem(clk, MemWrite, DataAdr, WriteData, MemReadData);
  
  // mux for switches:
  always_comb begin
        if (DataAdr == 32'hFF200040)
            ReadData = {22'b0, SW};   // Zero-extend 10-bit switches to 32-bit
        else
            ReadData = MemReadData;   // Default to Memory
  end

  always_ff @(posedge clk) begin
    if(reset) begin
      LEDR <= 10'b0;
      HEX3HEX0 <= 32'b0;
      HEX5HEX4 <= 16'b0;
    end
    else if (MemWrite) begin
      case(DataAdr)
        32'hFF200000:	LEDR <= WriteData[9:0];
        32'hFF200020:	HEX3HEX0 <= WriteData;
        32'hFF200030:	HEX5HEX4 <= WriteData[15:0];
      endcase
  	end
  end
      
  
endmodule

module riscvsingle(input logic clk, reset,
    output logic [31:0] PC,
    input logic [31:0] Instr,
    output logic MemWrite,
    output logic [31:0] ALUResult, WriteData,
    input logic [31:0] ReadData);

    logic ALUSrc, RegWrite, Jump, Zero, PCSrc;
    logic [1:0] ResultSrc, ImmSrc;
    logic [2:0] ALUControl;

    controller c(Instr[6:0], Instr[14:12], Instr[30], Zero,
                 ResultSrc, MemWrite, PCSrc,
                 ALUSrc, RegWrite, Jump,
                 ImmSrc, ALUControl);

    datapath dp(clk, reset, ResultSrc, PCSrc,
                ALUSrc, RegWrite,
                ImmSrc, ALUControl,
                Zero, PC, Instr,
                ALUResult, WriteData, ReadData);
endmodule

module controller(input logic [6:0] op,
    input logic [2:0] funct3,
    input logic funct7b5,
    input logic Zero,
    output logic [1:0] ResultSrc,
    output logic MemWrite,
    output logic PCSrc, ALUSrc,
    output logic RegWrite, Jump,
    output logic [1:0] ImmSrc,
    output logic [2:0] ALUControl);

    logic [1:0] ALUOp;
    logic Branch;

    maindec md(op, ResultSrc, MemWrite, Branch,
               ALUSrc, RegWrite, Jump, ImmSrc, ALUOp);

    aludec ad(op[5], funct3, funct7b5, ALUOp, ALUControl);

    assign PCSrc = Branch & Zero | Jump;
endmodule

module maindec(input logic [6:0] op,
    output logic [1:0] ResultSrc,
    output logic MemWrite,
    output logic Branch, ALUSrc,
    output logic RegWrite, Jump,
    output logic [1:0] ImmSrc,
    output logic [1:0] ALUOp);

    logic [10:0] controls;
    assign {RegWrite, ImmSrc, ALUSrc, MemWrite, ResultSrc, Branch, ALUOp, Jump} = controls;

    always_comb
        case(op)
            // RegWrite_ImmSrc_ALUSrc_MemWrite_ResultSrc_Branch_ALUOp_Jump
            7'b0000011: controls = 11'b1_00_1_0_01_0_00_0; // lw
            7'b0100011: controls = 11'b0_01_1_1_00_0_00_0; // sw
            7'b0110011: controls = 11'b1_xx_0_0_00_0_10_0; // R-type
            7'b1100011: controls = 11'b0_10_0_0_00_1_01_0; // beq
            7'b0010011: controls = 11'b1_00_1_0_00_0_10_0; // I-type ALU
            7'b1101111: controls = 11'b1_11_0_0_10_0_00_1; // jal
            default:    controls = 11'bx_xx_x_x_xx_x_xx_x; // ???
        endcase
endmodule

module aludec(input logic opb5,
    input logic [2:0] funct3,
    input logic funct7b5,
    input logic [1:0] ALUOp,
    output logic [2:0] ALUControl);

    logic RtypeSub;
    assign RtypeSub = funct7b5 & opb5; // TRUE for R-type subtract

    always_comb
        case(ALUOp)
            2'b00: ALUControl = 3'b000; // addition
            2'b01: ALUControl = 3'b001; // subtraction
            default: case(funct3) // R-type or I-type ALU
                3'b000: if (RtypeSub)
                            ALUControl = 3'b001; // sub
                        else
                            ALUControl = 3'b000; // add
                3'b010: ALUControl = 3'b101; // slt
                3'b110: ALUControl = 3'b011; // or, ori
                3'b111: ALUControl = 3'b010; // and, andi
                default: ALUControl = 3'bxxx;
            endcase
        endcase
endmodule

module datapath(input logic clk, reset,
    input logic [1:0] ResultSrc,
    input logic PCSrc, ALUSrc,
    input logic RegWrite,
    input logic [1:0] ImmSrc,
    input logic [2:0] ALUControl,
    output logic Zero,
    output logic [31:0] PC,
    input logic [31:0] Instr,
    output logic [31:0] ALUResult, WriteData,
    input logic [31:0] ReadData);

    logic [31:0] PCNext, PCPlus4, PCTarget;
    logic [31:0] ImmExt;
    logic [31:0] SrcA, SrcB;
    logic [31:0] Result;

    // next PC logic
    flopr #(32) pcreg(clk, reset, PCNext, PC);
    adder pcadd4(PC, 32'd4, PCPlus4);
    adder pcaddbranch(PC, ImmExt, PCTarget);
    mux2 #(32) pcmux(PCPlus4, PCTarget, PCSrc, PCNext);

    // register file logic
    regfile rf(clk, RegWrite, Instr[19:15], Instr[24:20], Instr[11:7], Result, SrcA, WriteData);
    extend ext(Instr[31:7], ImmSrc, ImmExt);

    // ALU logic
    mux2 #(32) srcbmux(WriteData, ImmExt, ALUSrc, SrcB);
    alu alu(SrcA, SrcB, ALUControl, ALUResult, Zero);
    mux3 #(32) resultmux(ALUResult, ReadData, PCPlus4, ResultSrc, Result);
endmodule

module extend(input logic [31:7] instr,
    input logic [1:0] immsrc,
    output logic [31:0] immext);

    always_comb
        case(immsrc)
            // I-type
            2'b00: immext = {{20{instr[31]}}, instr[31:20]};
            // S-type (stores)
            2'b01: immext = {{20{instr[31]}}, instr[31:25], instr[11:7]};
            // B-type (branches)
            2'b10: immext = {{20{instr[31]}}, instr[7], instr[30:25], instr[11:8], 1'b0};
            // J-type (jal)
            2'b11: immext = {{12{instr[31]}}, instr[19:12], instr[20], instr[30:21], 1'b0};
            default: immext = 32'bx; // undefined
        endcase
endmodule

module flopr #(parameter WIDTH = 8)
    (input logic clk, reset,
    input logic [WIDTH-1:0] d,
    output logic [WIDTH-1:0] q);

    always_ff @(posedge clk, posedge reset)
        if (reset) q <= 0;
        else q <= d;
endmodule

module flopenr #(parameter WIDTH = 8)
    (input logic clk, reset, en,
    input logic [WIDTH-1:0] d,
    output logic [WIDTH-1:0] q);

    always_ff @(posedge clk, posedge reset)
        if (reset) q <= 0;
        else if (en) q <= d;
endmodule

module mux2 #(parameter WIDTH = 8)
    (input logic [WIDTH-1:0] d0, d1,
    input logic s,
    output logic [WIDTH-1:0] y);

    assign y = s ? d1 : d0; // Fixed: was d1 : 0
endmodule

module mux3 #(parameter WIDTH = 8)
    (input logic [WIDTH-1:0] d0, d1, d2,
    input logic [1:0] s,
    output logic [WIDTH-1:0] y);

    assign y = s[1] ? d2 : (s[0] ? d1 : d0);
endmodule

module adder(input [31:0] a, b,
    output [31:0] y);
    assign y = a + b;
endmodule

module regfile(input logic clk,
    input logic we3,
    input logic [4:0] a1, a2, a3, // Fixed: was [5:0]
    input logic [31:0] wd3,
    output logic [31:0] rd1, rd2);

    logic [31:0] rf[31:0];

    // three ported register file
    // read two ports combinationally (A1/RD1, A2/RD2)
    // write third port on rising edge of clock (A3/WD3/WE3)
    // register 0 hardwired to 0
    always_ff @(posedge clk)
        if (we3) rf[a3] <= wd3;

    assign rd1 = (a1 != 0) ? rf[a1] : 0;
    assign rd2 = (a2 != 0) ? rf[a2] : 0;
endmodule

module alu(input logic [31:0] a, b,
    input logic [2:0] alucontrol,
    output logic [31:0] result,
    output logic zero);

    logic [31:0] condinvb, sum;
    logic v;
    logic isAddSub;

    assign condinvb = alucontrol[0] ? ~b : b;
    assign sum = a + condinvb + alucontrol[0];
    assign isAddSub = ~alucontrol[2] & ~alucontrol[1] | ~alucontrol[1] & alucontrol[0];

    always_comb
        case(alucontrol)
            3'b000: result = sum; // add
            3'b001: result = sum; // sub
            3'b010: result = a & b; // and
            3'b011: result = a | b; // or
            3'b100: result = a ^ b; // xor
            3'b101: result = sum[31] ^ v; // slt
            3'b110: result = a << b[4:0]; // sll
            3'b111: result = a >> b[4:0]; // srl
            default: result = 32'bx;
        endcase

    assign zero = (result == 32'b0);
    assign v = ~(alucontrol[0] ^ a[31] ^ b[31]) & (a[31] ^ sum[31]) & isAddSub;
endmodule

module imem(input logic [31:0] a,
    output logic [31:0] rd);

    logic [31:0] RAM[63:0];

    initial
      $readmemh("C:/Users/arvin/211/lab11/imem.txt", RAM);
    assign rd = RAM[a[31:2]]; // word aligned
endmodule

module dmem(input logic clk, we,
    input logic [31:0] a, wd,
    output logic [31:0] rd);

    logic [31:0] RAM[63:0]; // Fixed missing semicolon
	
  	initial
      $readmemh("C:/Users/arvin/211/lab11/dmem.txt", RAM);
  
    assign rd = RAM[a[31:2]]; // word aligned

    always_ff @(posedge clk)
        if (we) RAM[a[31:2]] <= wd;
endmodule